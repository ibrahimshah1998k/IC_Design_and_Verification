package my_testbench_pkg;
import uvm_pkg::*; 
`include "uvm_macros.svh"

`include "cc_seq_item.sv"
`include "cc_sequencer.sv"
`include "cc_sequence.sv"
`include "cc_driver.sv"
`include "cc_monitor.sv"
`include "cc_agent.sv"
`include "cc_scoreboard.sv"
`include "cc_env.sv"
`include "cc_base_test.sv"
endpackage
