package my_testbench_pkg;
import uvm_pkg::*; 
`include "uvm_macros.svh"

`include "mul_seq_item.sv"
`include "mul_sequencer.sv"
`include "mul_sequence.sv"
`include "mul_driver.sv"
`include "mul_monitor.sv"
`include "mul_agent.sv"
`include "mul_scoreboard.sv"
`include "mul_coverage.sv"
`include "mul_env.sv"
`include "mul_base_test.sv"
endpackage
