package my_testbench_pkg;
import uvm_pkg::*; 
`include "uvm_macros.svh"

`include "APB_seq_item.sv"
`include "APB_sequencer.sv"
`include "APB_sequence.sv"
`include "APB_driver.sv"
`include "APB_monitor.sv"
`include "APB_agent.sv"
`include "APB_scoreboard.sv"
`include "APB_env.sv"
`include "APB_base_test.sv"
endpackage
